package std_types;
	typedef logic bool;
	typedef logic [7:0] u8;
	typedef logic [15:0] u16;
	typedef logic [31:0] u32;
	typedef logic [63:0] u64;
	typedef logic [127:0] u128;
endpackage
